//写入管理模块，用于指挥Write Arbiter向SRAM中写入数据包

module write_manager();
    
endmodule 
