//用于寻找存储空间并维护链表

module space_finder();
    
endmodule 
