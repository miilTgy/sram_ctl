module arbiter_tb ();

    parameter arbiter_data_width = 256;
    reg ckl, rst;
    reg [arbiter_data_width-1:0] data_in;
    
endmodule