module arbiter_core_tb ();
    
endmodule