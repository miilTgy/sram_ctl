module fifo #(
  parameters
) (
  input data_in,
  output data_o
);
  
endmodule