module priority_decoder #(
    // parameters
) (
    // ports
);
    
endmodule