module cache_manager (
    input      clk,
    input      rst,
    
);
    
endmodule 
