module top (
    ports
);
    
endmodule