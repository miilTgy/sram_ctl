module ();

endmodule