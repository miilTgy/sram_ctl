module arbiter #(
    // parameters
) (
    // ports
);
    
endmodule