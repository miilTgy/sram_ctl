module ();
endmodule