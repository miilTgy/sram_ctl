module channel_selecter_tb ();
    parameter arbiter_data_width = 256;
    parameter num_of_ports = 16;
    reg clk, 
endmodule