module channel_selecter #(
    // parameters
) (
    // ports
);
    
endmodule