module arbiter_core (
    // ports
);
    
endmodule