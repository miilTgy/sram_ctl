//用于记录内存空间的链表，寻找内存可用空间和内存回收

module chain_manager();
    
endmodule 
