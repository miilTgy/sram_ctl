module ();
    parameter sg_data_width = 64;
    parameter sg_address_width = 12;
    parameter sg_des_width = 4;
    parameter sg_priority_width = 3;

endmodule