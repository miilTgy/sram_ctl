module fifo #(
  // parameters
  fifo_data_width = 256
) (
  // ports
  input data_in,
  output data_o
);
  
endmodule