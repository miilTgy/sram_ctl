module core_selecter_tb ();
endmodule