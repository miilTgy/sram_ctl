//用于记录内存空间状态的链表

module chain_recorder();
    
endmodule 
